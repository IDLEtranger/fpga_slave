`timescale 1ns / 1ps

module tb_pulse_statistic;